module stage2_tb; 






endmodule
